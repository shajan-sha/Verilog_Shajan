module HA_tb;
  
  reg a, b;
  wire s, c;
  
  
